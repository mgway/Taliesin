`timescale 1ns / 1ps

/* Taliesin Processor
 * 9/14/2013 - Version 1
 *
 * Description:
 * Work in progress
 * 
 */
 
module proc(
    );


endmodule
